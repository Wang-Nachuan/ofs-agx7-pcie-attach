//Copyright (C) 2021 Intel Corporation
//SPDX-License-Identifier: MIT
`ifndef TEST_TOP_PKG_NO_PMCI_SVH
`define TEST_TOP_PKG_NO_PMCI_SVH

    `include "test_pkg_no_pmci.svh"
    `include "test_long_pkg.svh"


`endif // TEST_TOP_PKG_NO_PMCI_SVH
